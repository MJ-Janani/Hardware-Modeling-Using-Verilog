module inverter(a,y);
input a;
output y;
not(y,a);
endmodule
